netcdf \20200101144000-ABOM-L3C_GHRSST-SSTskin-AHI_H08-1d_night-v02.0-fv02.0 {
dimensions:
	time = UNLIMITED ; // (1 currently)
	lat = 4500 ;
	lon = 6000 ;
variables:
	int time(time) ;
		time:_FillValue = -2147483647 ;
		time:long_name = "reference time of sst file" ;
		time:standard_name = "time" ;
		time:axis = "T" ;
		time:units = "seconds since 1981-01-01" ;
		time:comment = "A typical reference time for the data" ;
		time:calendar = "gregorian" ;
	float lat(lat) ;
		lat:_FillValue = 9.96921e+36f ;
		lat:long_name = "latitude" ;
		lat:standard_name = "latitude" ;
		lat:axis = "Y" ;
		lat:comment = "Latitudes for locating data" ;
		lat:valid_min = -90.f ;
		lat:valid_max = 90.f ;
		lat:units = "degrees_north" ;
	float lon(lon) ;
		lon:_FillValue = 9.96921e+36f ;
		lon:long_name = "longitude" ;
		lon:standard_name = "longitude" ;
		lon:axis = "X" ;
		lon:comment = "Longitudes for locating data" ;
		lon:valid_min = -180.f ;
		lon:valid_max = 360.f ;
		lon:units = "degrees_east" ;
	short sea_surface_temperature(time, lat, lon) ;
		sea_surface_temperature:_FillValue = -32768s ;
		sea_surface_temperature:add_offset = 289.59 ;
		sea_surface_temperature:scale_factor = 0.01 ;
		sea_surface_temperature:valid_min = -32765s ;
		sea_surface_temperature:valid_max = 32765s ;
		sea_surface_temperature:units = "kelvin" ;
		sea_surface_temperature:long_name = "sea surface skin temperature" ;
		sea_surface_temperature:standard_name = "sea_surface_skin_temperature" ;
		sea_surface_temperature:comment = "The skin temperature of the ocean at a depth of approximately 10 microns. SSTs are retrieved by using the Radiative Transfer Model (RTTOV12.3) and Bayesian cloud clearing method based on the ESA CCI SST code developed at the University of Reading" ;
		sea_surface_temperature:calendar = "Standard" ;
		sea_surface_temperature:coordinates = "time lat lon" ;
		sea_surface_temperature:grid_mapping = "crs" ;
	byte sses_bias(time, lat, lon) ;
		sses_bias:add_offset = 0. ;
		sses_bias:scale_factor = 0.00476172200395551 ;
		sses_bias:_FillValue = -128b ;
		sses_bias:valid_min = -127b ;
		sses_bias:valid_max = 127b ;
		sses_bias:clip_min = -0.604733932780346 ;
		sses_bias:clip_max = 0.504738558068635 ;
		sses_bias:units = "kelvin" ;
		sses_bias:long_name = "SSES bias estimate" ;
		sses_bias:comment = "Bias estimate derived from L2P bias,following the method described in http://imos.org.au/fileadmin/user_upload/shared/SRS/SST/GHRSST-DOC-basic-v1.0r1.pdf. Subtracting sses_bias from sea_surface_temperature produces a more accurate skin SST estimate" ;
		sses_bias:coordinates = "time lat lon" ;
		sses_bias:grid_mapping = "crs" ;
	byte sses_standard_deviation(time, lat, lon) ;
		sses_standard_deviation:add_offset = 0.805315375788983 ;
		sses_standard_deviation:scale_factor = 0.00241112387960773 ;
		sses_standard_deviation:_FillValue = -128b ;
		sses_standard_deviation:valid_min = -127b ;
		sses_standard_deviation:valid_max = 127b ;
		sses_standard_deviation:clip_min = 0.5 ;
		sses_standard_deviation:clip_max = 1.11242064317261 ;
		sses_standard_deviation:units = "kelvin" ;
		sses_standard_deviation:long_name = "SSES standard deviation estimate" ;
		sses_standard_deviation:comment = "Standard deviation estimate derived from L2P standard deviation, following the method described in http://imos.org.au/fileadmin/user_upload/shared/SRS/SST/GHRSST-DOC-basic-v1.0r1.pdf." ;
		sses_standard_deviation:coordinates = "time lat lon" ;
		sses_standard_deviation:grid_mapping = "crs" ;
	byte quality_level(time, lat, lon) ;
		quality_level:add_offset = 0. ;
		quality_level:scale_factor = 1. ;
		quality_level:_FillValue = -128b ;
		quality_level:valid_min = -127b ;
		quality_level:valid_max = 127b ;
		quality_level:long_name = "quality level of SST pixel" ;
		quality_level:comment = "These are the overall quality indicators and are used for all GHRSST SSTs. Refer Merchant et al., 2019 (https://doi.org/10.1038/s41597-019-0236-x) for more details for logic and threshold for assigning pixel quality level with use of Bayesian cloud clearing method. For validation applications, please consider quality_level greater than or equal 4 with bias correction. For operational applications, please consider quality_level greater than or equal 4 with bias correction. For qualitative applications, please consider quality_level greater than or equal 3 with or without bias correction." ;
		quality_level:flag_meanings = "no_data bad_data worst_quality low_quality acceptable_quality best_quality" ;
		quality_level:coordinates = "time lat lon" ;
		quality_level:grid_mapping = "crs" ;
		quality_level:flag_values = 0b, 1b, 2b, 3b, 4b, 5b ;
	short sst_dtime(time, lat, lon) ;
		sst_dtime:_FillValue = -32768s ;
		sst_dtime:add_offset = -300. ;
		sst_dtime:scale_factor = 1. ;
		sst_dtime:valid_min = -32765s ;
		sst_dtime:valid_max = 32765s ;
		sst_dtime:units = "second" ;
		sst_dtime:long_name = "time difference from reference time" ;
		sst_dtime:comment = "time plus sst_dtime gives seconds after 00:00:00 UTC January 1, 1981." ;
		sst_dtime:coordinates = "time lat lon" ;
		sst_dtime:grid_mapping = "crs" ;
	byte dt_analysis(time, lat, lon) ;
		dt_analysis:add_offset = 0. ;
		dt_analysis:scale_factor = 0.1 ;
		dt_analysis:_FillValue = -128b ;
		dt_analysis:valid_min = -127b ;
		dt_analysis:valid_max = 127b ;
		dt_analysis:units = "Kelvin" ;
		dt_analysis:long_name = "deviation from last SST analysis" ;
		dt_analysis:comment = "The difference between this SST and the previous day\'s L4 Foundation SST." ;
		dt_analysis:source = "ABOM-L4LRfnd-GLOB-GAMSSA_28km" ;
		dt_analysis:coordinates = "time lat lon" ;
		dt_analysis:grid_mapping = "crs" ;
	short l2p_flags(time, lat, lon) ;
		l2p_flags:_FillValue = -32768s ;
		l2p_flags:valid_min = -32765s ;
		l2p_flags:valid_max = 32765s ;
		l2p_flags:long_name = "L2P flags" ;
		l2p_flags:comment = "These flags are important to properly use the data.  Data not flagged as microwave are sourced from an infrared sensor. The lake and river flags are currently not set, but defined in GDS2.0r4. The terminator flag indicates that the sun is near the horizon. The analysis flag indicates high difference from analysis temperatures (differences greater than Analysis Limit). The lowwind flag indicates regions of low wind speed (typically less than the low Wind Limit) per NWP model. The highwind flag indicates regions of high wind speed (typically greater than the high Wind Limit) per NWP model. Other flags may be populated and are for internal use and the definitions may change, so should not be relied on. Use flag_meanings to confirm the flag assignment that can be relied on. Flags greater than 64 only apply to non-land pixels." ;
		l2p_flags:coordinates = "time lat lon" ;
		l2p_flags:grid_mapping = "crs" ;
		l2p_flags:flag_masks = 1s, 2s, 4s, 8s, 16s, 32s, 64s, 128s, 256s, 512s, 1024s, 2048s, 4096s, 8192s, 16384s ;
		l2p_flags:flag_meanings = "microwave land ice lake river reserved reserved analysis lowwind highwind night terminator reserved reserved reserved" ;
	byte sses_count(time, lat, lon) ;
		sses_count:add_offset = 14.0919070602216 ;
		sses_count:scale_factor = 0.10286063547607 ;
		sses_count:_FillValue = -128b ;
		sses_count:valid_min = -127b ;
		sses_count:valid_max = 127b ;
		sses_count:clip_min = 0.992141608467754 ;
		sses_count:clip_max = 27.1185372981186 ;
		sses_count:units = "count" ;
		sses_count:long_name = "SSES count" ;
		sses_count:comment = "Weighted representative number of swath pixels, per https://imos.org.au/facilities/srs/sstproducts/sstdata0/sstdata-ghrsstfilefields. EXPERIMENTAL_FIELD" ;
		sses_count:coordinates = "time lat lon" ;
		sses_count:grid_mapping = "crs" ;
	byte wind_speed(time, lat, lon) ;
		wind_speed:add_offset = 8.7125486893654 ;
		wind_speed:scale_factor = 0.0686027455855543 ;
		wind_speed:_FillValue = -128b ;
		wind_speed:valid_min = -127b ;
		wind_speed:valid_max = 127b ;
		wind_speed:clip_min = 0. ;
		wind_speed:clip_max = 17.4249601732396 ;
		wind_speed:long_name = "wind_speed" ;
		wind_speed:standard_name = "wind_speed" ;
		wind_speed:comment = "Typically represent surface winds (10 meters above the sea surface)." ;
		wind_speed:source = "ACCESSG-ABOM-Forecast-WSP" ;
		wind_speed:coordinates = "time lat lon" ;
		wind_speed:grid_mapping = "crs" ;
		wind_speed:units = "m s-1" ;
	byte satellite_zenith_angle(time, lat, lon) ;
		satellite_zenith_angle:add_offset = 35.0459746431039 ;
		satellite_zenith_angle:scale_factor = 0.275952556244913 ;
		satellite_zenith_angle:_FillValue = -128b ;
		satellite_zenith_angle:valid_min = -127b ;
		satellite_zenith_angle:valid_max = 127b ;
		satellite_zenith_angle:clip_min = 0. ;
		satellite_zenith_angle:clip_max = 70.0913973810954 ;
		satellite_zenith_angle:units = "angular_degree" ;
		satellite_zenith_angle:long_name = "satellite_zenith angle" ;
		satellite_zenith_angle:comment = "The satellite zenith angle at the time of the SST observations" ;
		satellite_zenith_angle:coordinates = "time lat lon" ;
		satellite_zenith_angle:grid_mapping = "crs" ;
	byte sea_ice_fraction(time, lat, lon) ;
		sea_ice_fraction:add_offset = 0. ;
		sea_ice_fraction:scale_factor = 1. ;
		sea_ice_fraction:_FillValue = -128b ;
		sea_ice_fraction:valid_min = -127b ;
		sea_ice_fraction:valid_max = 127b ;
		sea_ice_fraction:units = "1" ;
		sea_ice_fraction:long_name = "sea_ice_fraction" ;
		sea_ice_fraction:standard_name = "sea_ice_area_fraction" ;
		sea_ice_fraction:comment = "Fractional sea ice cover (unitless) derived from near real-time UKMO OSTIA Daily 0.05 degree L4, an optimal interpolation of the operational near real-time EUMETSAT OSI-SAF SSMIS daily 10 km Level 3 sea ice concentration fields (Good et al., 2020, Remote Sensing, https://dx.doi.org/10.3390/rs12040720)." ;
		sea_ice_fraction:source = "OSTIA-UKMO-L4-GLOB-v2.0" ;
		sea_ice_fraction:coordinates = "time lat lon" ;
		sea_ice_fraction:grid_mapping = "crs" ;
	int crs ;
		crs:long_name = "coordinate reference system" ;
		crs:grid_mapping_name = "latitude_longitude" ;
		crs:semi_major_axis = 6379137.f ;
		crs:inverse_flattening = 298.257223563 ;
		crs:epsg_code = "EPSG:4326" ;

// global attributes:
		:id = "AHI_H08-ABOM-L3C-v02.0" ;
		:Conventions = "CF-1.6" ;
		:title = "Nighttime gridded single-sensor multiple-swath Australian region Himawari-8 AHI SST" ;
		:summary = "Skin sea surface temperature retrievals from the AHI sensor on the Himawari-8 satellite, regridded IMOS L3C-01day night SST on native grid to 0.02 degree rectangular grid over the Australian domain, produced by the Australian Bureau of Meteorology in collaboration with University of Reading" ;
		:references = "https://www.foo.org.au/wp-content/uploads/2021/11/Govekar_FOO_2021.pdf, http://imos.org.au/sstproducts.html, https://doi.org/10.1038/s41597-019-0236-x, http://imos.org.au/fileadmin/user_upload/shared/SRS/SST/GHRSST-DOC-basic-v1.0r1.pdf, https://zenodo.org/record/4700466" ;
		:institution = "ABOM" ;
		:comment = "Multi swath AHI_H08  SSTskin retrievals obtained from regridding IMOS Himawari-8 L3C-01day night file on native grid, produced by the Australian Bureau of Meteorology. This is gridded SST defined on 0.02 degree rectangular grid over the Australian domain for the night (before dawn). SSTs were retrieved by using the Radiative Transfer Model (RTTOV12.3) and Bayesian cloud clearing method based on the ESA CCI SST code developed at the University of Reading." ;
		:license = "GHRSST protocol describes data use as free and open" ;
		:naming_authority = "org.ghrsst" ;
		:product_version = "2.0" ;
		:uuid = "ea7c053e-1589-4259-a7ab-805e433bb262" ;
		:gds_version_id = "2.0r5" ;
		:netcdf_version_id = "4.6." ;
		:spatial_resolution = "0.02 deg" ;
		:platform = "Himawari-8" ;
		:sensor = "AHI" ;
		:Metadata_Conventions = "Unidata Observation Dataset v1.0" ;
		:Metadata_Link = "TBA" ;
		:keywords = "Oceans > Ocean Temperature > Sea Surface Temperature" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords" ;
		:standard_name_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Convention" ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_units = "degrees_east" ;
		:geospatial_lat_resolution = 0.02f ;
		:geospatial_lon_resolution = 0.02f ;
		:notes = "quality=archive" ;
		:history = "sst_source=AHI_H08-ABOM-L3C-night_Geos141-v02.0,wind_source=ACCESSG-ABOM-Analysis-WSP,ACCESSG-ABOM-Forecast-WSP,analysis_source=ABOM-L4LRfnd-GLOB-GAMSSA_28km,analysis_file=20191231-ABOM-L4LRfnd-GLOB-v01-fv01.nc,ice_source=OSTIA-UKMO-L4-GLOB-v2.0,ice_file=20200101120000-UKMO-L4_GHRSST-SSTfnd-OSTIA-GLOB-v02.0-fv02.0.nc,NoWindForecast=0,NoIce=0,qssesscale=-0.143,qsseszero=0.25,qssesdone=0,quality=archive" ;
		:acknowledgment = "Any use of these data requires the following acknowledgment:\"AHI SSTskin retrieval produced by the Australian Bureau of Meteorology, in collaboration with University of Reading as a contribution to the Integrated Marine Observing System (IMOS) - IMOS is enabled by the National Collaborative Research Infrastructure (NCRIS). The imagery data are acquired from the Himawari-8 spacecraft by the Japan Aerospace Exploration Agency." ;
		:creator_name = "Australian Bureau of Meteorology" ;
		:creator_email = "ghrsst@bom.gov.au" ;
		:creator_url = "http://www.bom.gov.au" ;
		:project = "Group for High Resolution Sea Surface Temperature" ;
		:publisher_name = "The GHRSST Project Office" ;
		:publisher_email = "gpa@ghrsst.org" ;
		:publisher_url = "http://www.ghrsst.org" ;
		:processing_level = "L3C" ;
		:cdm_data_type = "Grid" ;
		:date_created = "20220726T222829Z" ;
		:start_time = "20200101T034000Z" ;
		:time_coverage_start = "20200101T034000Z" ;
		:stop_time = "20200102T034000Z" ;
		:time_coverage_end = "20200102T034000Z" ;
		:file_quality_level = 3 ;
		:northernmost_latitude = "19.99f" ;
		:southernmost_latitude = "-69.99f" ;
		:easternmost_longitude = "-170.01f" ;
		:westernmost_longitude = "70.01f" ;
		:source = "wind_source=ACCESSG-ABOM-Forecast-WSP,analysis_source=ABOM-L4LRfnd-GLOB-GAMSSA_28km,ice_source=OSTIA-UKMO-L4-GLOB-v2.0,l2_source=AHI_H08-ABOM-L2P-v02.0" ;
}
